---------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- Course: University of Victoria
-- Engineer: Jake Friesen, Matthew Ebert, Samuel Pacheo 
-- 
-- Create Date: 2023-Mar-09

-- Module Name: Write_Back_Stage - Behavioral
-- Project Name: 16bitCPU
-- Target Devices: Artix7
-- Description: 
-- 
-- Dependencies: 
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library work;
use work.Constant_Package.all;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;


entity Memory_Stage is
    Port ( Result_MEM_in : in STD_LOGIC_VECTOR (15 downto 0);
           IR_MEM_in : in STD_LOGIC_VECTOR (15 downto 0);
           clk, rst : in STD_LOGIC;
           branch_flush : in std_logic;
           ram_wren_A: out std_logic;
           ram_en_A: out std_logic;
           ram_wrdata_A: out STD_LOGIC_VECTOR (15 downto 0);
           ram_addr_A: out std_logic_vector (15 downto 0);
           ram_data_A: in std_logic_vector (15 downto 0);
           memdata_MEM_out : out STD_LOGIC_VECTOR (15 downto 0);
           Result_MEM_out : out STD_LOGIC_VECTOR (15 downto 0);
           IR_MEM_out : out STD_LOGIC_VECTOR (15 downto 0);
           vdata_MEM_in, A_MEM_in, B_MEM_in : in STD_LOGIC_VECTOR (15 downto 0);
           vdata_MEM_out : out STD_LOGIC_VECTOR (15 downto 0));
end Memory_Stage;

architecture Behavioral of Memory_Stage is
    signal IR, ALU, Overflow, ram_output : std_logic_vector (15 downto 0);

begin
    --Latch Process
    process(clk)
    begin
        if(rst = '1') then
        --Reset
            IR_MEM_out <= (others=>'0');
            vdata_MEM_out <= (others=>'0');
            Result_MEM_out <= (others=>'0');
            memdata_MEM_out <= (others=>'0');  
        end if;    
        if(clk'event and clk = '1') then
        --Latch Incoming signals
            if(branch_flush = '1') then
            --Internal Branch set, clear the incoming buffer
                IR <= (others=>'0');
                ALU <= (others=>'0');
                Overflow <= (others=>'0');
            else
                IR <= IR_MEM_in;
                ALU <= Result_MEM_in;
                Overflow <= vdata_MEM_in;
            end if;
        end if;
        if(clk'event and clk = '0') then
        --Latch Outgoing signals
            vdata_MEM_out <= Overflow;
            IR_MEM_out <= IR;
            Result_MEM_out <= ALU;
            
            if(IR(15 downto 9) = mov_op or IR(15 downto 9) = out_op) then
                memdata_MEM_out <= A_MEM_in;
            else
                memdata_MEM_out <= ram_data_A;
            end if;  
                
        end if;
    end process;

    --RAM Access
    with IR_MEM_in(15 downto 9) Select
        ram_wren_A <=   '1' when store_op | push_op, --STR (17), PUSH (96)
                    '0' when others;  
                    
    with IR_MEM_in(15 downto 9) Select
         ram_en_A <=  '1' when store_op | load_op | push_op | pop_op,
                     '0' when others;  
    
    ram_addr_A <= A_MEM_in(15 downto 0);
    ram_wrdata_A <=  B_MEM_in;
    
end Behavioral;